`define DELAY 20
module alu_testbench(); 
reg [31:0]A, B;
reg carry_in;
reg [2:0] S;
wire [31:0]result;


alu g0(A, B,S,carry_in,result);



initial begin
A = 32'b0000_0000_0000_0000_0000_0000_0000_1101; B = 32'b0000_0000_0000_0000_0000_0000_0000_1001; carry_in = 1'b0; S = 3'b000;
#`DELAY;
A = 32'b0000_0000_0000_0000_0000_0000_0000_1011; B = 32'b0000_0000_0000_0000_0000_0000_0000_1110; carry_in = 1'b0; S = 3'b001;
#`DELAY;
A = 32'b0000_0000_0000_0000_0000_0000_0000_1111; B = 32'b0000_0000_0000_0000_0000_0000_0000_1010; carry_in = 1'b0; S = 3'b010;
#`DELAY;
A = 32'b0000_0000_0000_0000_0000_0000_0000_0001; B = 32'b0000_0000_0000_0000_0000_0000_0000_1101; carry_in = 1'b0; S = 3'b011;
#`DELAY;
A = 32'b0000_0000_0000_0000_0000_0000_0000_1011; B = 32'b0000_0000_0000_0000_0000_0000_0000_0110; carry_in = 1'b0; S = 3'b100;
#`DELAY;
A = 32'b0000_0000_0000_0000_0000_0000_0000_0011; B = 32'b0000_0000_0000_0000_0000_0000_0000_0011; carry_in = 1'b0; S = 3'b101;
#`DELAY;
A = 32'b0000_0000_0000_0000_0000_0000_0000_0100; B = 32'b0000_0000_0000_0000_0000_0000_0000_1111; carry_in = 1'b0; S = 3'b110;
#`DELAY;
A = 32'b0000_0000_0000_0000_0000_0000_0000_1001; B = 32'b0000_0000_0000_0000_0000_0000_0000_0100; carry_in = 1'b0; S = 3'b111;
#`DELAY;


end
 
 
initial
begin
$monitor("time = %2d, a =%32b, b=%32b , S=%3b, result=%32b", $time, A, B , S, result);
end
 
endmodule